interface fa_intf;
  logic a;
  logic b;
  logic cin;
  logic sum;
  logic cout;
endinterface
